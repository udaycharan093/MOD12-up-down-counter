/********************************************************************************************

Copyright 2019 - Maven Silicon Softech Pvt Ltd.  
www.maven-silicon.com

All Rights Reserved.

This source code is an unpublished work belongs to Maven Silicon Softech Pvt Ltd.
It is not to be shared with or used by any third parties who have not enrolled for our paid 
training courses or received any written authorization from Maven Silicon.

Filename       :  ram_read_mon.sv   

Description    :  Monitor class for dual port ram_testbench

Author Name    :  Putta Satish

Support e-mail :  techsupport_vm@maven-silicon.com 

Version        :  1.0

Date           :  02/06/2020

***********************************************************************************************/
//In class ram_read_mon

class mod_read_mon;

   //Instantiate virtual interface instance rd_mon_if of type ram_if with RD_MON_MP modport
   virtual mod_if.RD_MON_MP rd_mon_if;

   //Declare three handles 'rddata', 'data2rm' and 'data2sb' of class type ram_trans
   mod_trans rddata, data2sb;
// mod_trans data2rm;

   //Declare two mailboxes 'mon2rm' and 'mon2sb' parameterized by type ram_trans
// mailbox #(mod_trans) mon2rm;
   mailbox #(mod_trans) mon2sb;
   
   //In constructor
   //Pass the following as the input arguments  
   //virtual interface 
   //mailbox handles 'mon2rm' and 'mon2sb' parameterized by ram_trans   
   //make the connections and allocate memory for 'rddata'

   function new(virtual mod_if.RD_MON_MP rd_mon_if,
                mailbox #(mod_trans) mon2sb);
      this.rd_mon_if = rd_mon_if;
//      this.mon2rm    = mon2rm;
      this.mon2sb    = mon2sb;
      this.rddata    = new;
   endfunction: new


   virtual task monitor();
      @(rd_mon_if.rd_mon_cb);
      begin
         rddata.d_out = rd_mon_if.rd_mon_cb.d_out;
         //call the display of the ram_trans to display the monitor data
        // rddata.display("DATA FROM READ MONITOR");    
      end
   endtask: monitor
   
   
   //In virtual task start       
   virtual task start();
      //within fork-join_none
      //In forever loop
      fork
         forever
            begin
               //Call the monitor task
               //Understand the provided monitor task 
               //Monitor task samples the interface signals 
               //according to the protocol and convert to transaction items 
               monitor(); 

               //Shallow copy rddata to data2sb;
               //Shallow copy rddata to data2rm;
               data2sb = new rddata;
//	$display("%0d",data2sb.d_out);

//               data2rm = new rddata;
               //Put the transaction item into two mailboxes mon2rm and mon2sb
//               mon2rm.put(data2rm);
               mon2sb.put(data2sb);
			data2sb.display("Data From Read Monitor");
            end
      join_none
   endtask: start

endclass: mod_read_mon
